module tb ;

initial begin
$display("hell0");
end 
endmodule