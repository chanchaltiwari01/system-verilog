module print();
rag a = 1 , b=0 ;
initial begin
$display("a:%0d,b:%0d",a,b);
end 
initial begin
    $display("first change ");
end
endmodule 
