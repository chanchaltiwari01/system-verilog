module 
endmodule 
